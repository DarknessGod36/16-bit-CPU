module MiniProject (
    
);
    
endmodule